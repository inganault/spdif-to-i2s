module main (
  input wire clk, // 12.0MHz
  input wire pause,
  output reg drive_p
);


endmodule